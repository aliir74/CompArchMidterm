library verilog;
use verilog.vl_types.all;
entity myClock is
end myClock;
