module MainMem;  

reg [15:0] mem [0:8191];

endmodule
