library verilog;
use verilog.vl_types.all;
entity Cache_tb is
end Cache_tb;
