library verilog;
use verilog.vl_types.all;
entity Clock is
end Clock;
